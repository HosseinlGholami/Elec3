** Profile: "SCHEMATIC1-spaze2"  [ E:\AZ\2\paze2-schematic1-spaze2.sim ] 

** Creating circuit file "paze2-schematic1-spaze2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 30 7meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze2-SCHEMATIC1.net" 


.END
