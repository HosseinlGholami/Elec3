** Profile: "SCHEMATIC1-spaze8"  [ E:\AZ\8\paze8-schematic1-spaze8.sim ] 

** Creating circuit file "paze8-schematic1-spaze8.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze8-SCHEMATIC1.net" 


.END
