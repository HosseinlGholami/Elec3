** Profile: "SCHEMATIC1-spaze8-2"  [ E:\AZ\8\paze8-1-SCHEMATIC1-spaze8-2.sim ] 

** Creating circuit file "paze8-1-SCHEMATIC1-spaze8-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1 1 5000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze8-1-SCHEMATIC1.net" 


.END
