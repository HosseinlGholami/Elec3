** Profile: "SCHEMATIC1-spaze6"  [ E:\AZ\6\paze6-2-schematic1-spaze6.sim ] 

** Creating circuit file "paze6-2-schematic1-spaze6.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 100n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze6-2-SCHEMATIC1.net" 


.END
