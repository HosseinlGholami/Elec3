** Profile: "SCHEMATIC1-spaze3"  [ E:\AZ\3\paze3-schematic1-spaze3.sim ] 

** Creating circuit file "paze3-schematic1-spaze3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 10000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze3-SCHEMATIC1.net" 


.END
