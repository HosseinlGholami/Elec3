** Profile: "SCHEMATIC1-spaze7"  [ E:\AZ\7\paze7-schematic1-spaze7.sim ] 

** Creating circuit file "paze7-schematic1-spaze7.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paze7-SCHEMATIC1.net" 


.END
