** Profile: "SCHEMATIC1-spaze1"  [ E:\AZ\1\paz1-schematic1-spaze1.sim ] 

** Creating circuit file "paz1-schematic1-spaze1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 3 8meg
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\paz1-SCHEMATIC1.net" 


.END
